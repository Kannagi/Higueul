[build-menu]
FT_00_LB=
FT_00_CM=bash compile.sh
FT_00_WD=
EX_00_LB=_Exécuter
EX_00_CM=gtkwave prg.vcd
EX_00_WD=
